module test;
  reg [1:0] pattin;
  wire a, b;
  wire [1:0] o, pattout;
  reg [10*8:0] patFile, fltFile, rptFile;
  
  assign {a, b} = pattin;
  assign pattout = o;
  gate g1(o, a, b);
  initial
  begin   
    patFile = "pat.txt";
    fltFile = "fault.txt";
    rptFile = "fault.rpt";
    $faultEnumerate(fltFile);
    $generatePatterns(pattin, pattout, fltFile, patFile, rptFile);
  end                     
endmodule                 

module gate (
o,
a,
b
);
input  a;
input  b;
output [1:0] o;
// concat starts line no 4
buf (o[0], a);
buf (o[1], b);
// concat ends line no 4
endmodule
